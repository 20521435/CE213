`timescale 10ns/10ps
module tb_datapath ();
  reg CLK, regDst, regWrite, ALUSrc, ALUcontrol, memWrite, memRead, memtoReg;
  reg [31:0] INST;
  wire [31:0] regW, addr;
  wire isZero;
  datapath u1 (CLK, INST, regDst, regWrite, ALUSrc, ALUcontrol, memWrite, memRead, memtoReg, regW, isZero, addr);
  
  initial begin 
    CLK = 0; 
    INST = 32'b00000010010100111000100000100000;
    #10 //add $1, $2, $3
    regDst = 1; 
    regWrite = 0; 
    ALUSrc = 0; 
    ALUcontrol = 4'b0010; 
    memWrite = 0; 
    memRead = 0; 
    memtoReg = 0;
    #20
    regWrite = 1; 
    $monitor ("regW: %d", regW);
  end 
  always #10 CLK = ~CLK;
endmodule