library verilog;
use verilog.vl_types.all;
entity tb_process is
end tb_process;
